`timescale 1ns / 1ps

package spmv_pkg;


endpackage : spmv_pkg
