`timescale 1ns / 1ps

import spmv_pkg::*;

module spmv_network_op #(
) (
    input wire clk,
    input wire rst_n
);

endmodule

