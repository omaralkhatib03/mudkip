`timescale 1 ps/1 ps

module top#(

  ) (
    input wire                          clk,
    input wire                          rst_n,

  );


endmodule
