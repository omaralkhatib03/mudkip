`timescale 1ns / 1ps

package spmv_pkg;

typedef logic [63:0] long;


endpackage : spmv_pkg
