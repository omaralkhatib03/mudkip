`timescale 1ns/1ps

module attach_start_to_stream (
  input clk,
  input rst_n,

  axi_stream_if.slave in,
  axi_stream_if.master out
);


endmodule
