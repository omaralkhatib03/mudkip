`timescale 1 ns/1 ps

module top #(
) (
);

endmodule
