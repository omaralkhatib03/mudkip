`timescale 1ns / 1ps

module spmv_network_op_tb #(
) (
    input wire clk,
    input wire rst_n

);

endmodule
